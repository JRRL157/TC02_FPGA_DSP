`ifndef DP_RAM_CONTROLLER_DEFINES_V
`define DP_RAM_CONTROLLER_DEFINES_V

typedef enum logic [3:0] {
   ST_IDLE_RAM_CONTROLLER = 4'b000, 
	ST_WAIT_READ = 4'b0111,
	ST_READ_INPUT = 4'b0001, 
	ST_WAIT_OPERATION = 4'b0010,
	ST_WRITE_OUTPUT = 4'b0011,
	ST_WAIT_FINISH = 4'b1000,
	ST_SET_FINISH = 4'b0100,
	ST_WAIT_SHUTDOWN = 4'b0101,
	ST_CLEAR = 4'b0110
} dp_ram_controller_states_t;

`endif